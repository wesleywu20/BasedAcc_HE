module top;

    multiplier_itf itf();
    testbench tb (.*);
endmodule : top
