package rv32i_types;
// Mux types are in their own packages to prevent identiier collisions
// e.g. pcmux::pc_plus4 and regfilemux::pc_plus4 are seperate identifiers
// for seperate enumerated types
import pcmux::*;
import marmux::*;
import cmpmux::*;
import alumux::*;
import regfilemux::*;

typedef logic [31:0] rv32i_word;
typedef logic [4:0] rv32i_reg;
typedef logic [3:0] rv32i_mem_wmask;

typedef enum bit [6:0] {
    op_lui   = 7'b0110111, //load upper immediate (U type)
    op_auipc = 7'b0010111, //add upper immediate PC (U type)
    op_jal   = 7'b1101111, //jump and link (J type)
    op_jalr  = 7'b1100111, //jump and link register (I type)
    op_br    = 7'b1100011, //branch (B type)
    op_load  = 7'b0000011, //load (I type)
    op_store = 7'b0100011, //store (S type)
    op_imm   = 7'b0010011, //arith ops with register/immediate operands (I type)
    op_reg   = 7'b0110011, //arith ops with register operands (R type)
    op_csr   = 7'b1110011,  //control and status register (I type)
	op_accel = 7'b1111111
} rv32i_opcode;


typedef struct{
	bit [4:0] reg_id;
	bit [31:0] data;
}command_buffer;

typedef enum bit [2:0] {
    beq  = 3'b000,
    bne  = 3'b001,
    blt  = 3'b100,
    bge  = 3'b101,
    bltu = 3'b110,
    bgeu = 3'b111
} branch_funct3_t;

typedef enum bit [2:0] {
    lb  = 3'b000,
    lh  = 3'b001,
    lw  = 3'b010,
    lbu = 3'b100,
    lhu = 3'b101
} load_funct3_t;

typedef enum bit [2:0] {
    sb = 3'b000,
    sh = 3'b001,
    sw = 3'b010
} store_funct3_t;

typedef enum bit [2:0] {
    add  = 3'b000, //check bit30 for sub if op_reg opcode
    sll  = 3'b001,
    slt  = 3'b010,
    sltu = 3'b011,
    axor = 3'b100,
    sr   = 3'b101, //check bit30 for logical/arithmetic
    aor  = 3'b110,
    aand = 3'b111
} arith_funct3_t;

typedef enum bit [3:0] {
    alu_add = 4'b000,
    alu_sll = 4'b001,
    alu_sra = 4'b010,
    alu_sub = 4'b011,
    alu_xor = 4'b100,
    alu_srl = 4'b101,
    alu_or  = 4'b110,
    alu_and = 4'b111,
    alu_sltu = 4'b1000,
    alu_slt = 4'b1001
} alu_ops;


//Struct of the decoded instruction 
typedef struct  packed{
    bit [2:0] funct3;
    bit [6:0] funct7;
    rv32i_opcode opcode;
    bit [31:0] i_imm;
    bit [31:0] s_imm;
    bit [31:0] b_imm;
    bit [31:0] u_imm;
    bit [31:0] j_imm;
    bit [4:0] rs1;
    bit [4:0] rs2;
    bit [4:0] rd;
    bit [31:0] pc;
    bit [31:0] instruction;
	bit [2:0] branch_id;
} instr_struct;

parameter int width_p = $bits(instr_struct);
typedef logic [width_p-1:0] word_t;
// FIFO's don't use shift registers, rather, they use pointers
// which address to the "read" (dequeue) and "write" (enqueue)
// ports of the FIFO's memory
parameter int ptr_width_p = 2;

// Why is the ptr type a bit longer than the "ptr_width"? 
// Make sure you can answer this question by the end of the semester
typedef logic [ptr_width_p:0] ptr_t;

// The number of words stored in the FIFO
parameter int cap_p = 1 << ptr_width_p;

endpackage : rv32i_types

