module top;

    polymult_itf itf();
    polymult_tb tb (.*);

endmodule