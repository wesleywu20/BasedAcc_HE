`ifndef mult_constants
`define mult_constants

/* comment out whichever one based on which one you want to test */
// `define test_full_mult
// `define test_half_mult
`define test_param_mult

`define HALF_PROD_MASK 64'hFFFFFFFFFFFFFFFF

`endif