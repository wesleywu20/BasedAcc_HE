// Import parameters from file
`include "he_params.sv"

`resetall
